module and1(y,a,b);
    output y;
    input a,b;
    and g1(y,a,b);
endmodule